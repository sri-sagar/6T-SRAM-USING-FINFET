*sram cmos
*drain gate source bulk type

M1 qb q vdd vdd pmos w=120n l=45n
M2 q qb vdd vdd pmos w=120n l=45n
M3 q qb gnd gnd nmos w=120n l=45n
M4 qb q gnd gnd nmos w=120n l=45n
M5 qb wl blb gnd nmos w=120n l=45n
M6 q wl bl gnd nmos w=120n l=45n


* vwl word line WL
vwl wl 0 1

* vbl bit line BL
vbl bl 0 pulse(0 1 0.01n 1p 1p 10n 20n)

* vblb bit line bar BLB
vblb blb 0 pulse(1 0 0.01n 1p 1p 10n 20n)

*VDD
vdd vdd 0 1


.param supply=1.0
*transient analysis
.tran 1n 60n start=0
*.measure tran averagepower AVG POWER from 1n to 60n
.measure tran SupplyCurrent avg i(vdd) from 1n to 60n
.measure tran  DynamicPower PARAM='-SupplyCurrent*supply'
.print tran TotalPower total power from 1n to 60n


* PTM 32nm

.model  nmos  nmos  level = 54

+version = 4.0          binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 1          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0          

+tnom    = 27           toxe    = 1.4e-009     toxp    = 0.8e-009    toxm    = 1.4e-009   
+dtox    = 0.6e-9      epsrox  = 3.9          wint    = 0            lint    = 8.5e-009   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 1.4e-009   

+vth0    = 0.42252      k1      = 0.5          k2      = 0.05            k3      = 0          
+k3b     = 0            w0      = 0.0e-006     dvt0    = 1            dvt1    = 0.95       
+dvt2    = 0            dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 0.36         minv    = 0.0          voffl   = 0            dvtp0   = 0    
+dvtp1   = 0.0          lpe0    = 0            lpeb    = 0            xj      = 5e-008     
+ngate   = 5e+020       ndep    = 4.1e+018     nsd     = 2e+020       phin    = 0         
+cdsc    = 0.07         cdscb   = 0            cdscd   = 0.02          cit     = 0          
+voff    = -0.09        nfactor = 1.5          eta0    = 0.035         etab    = 0          
+vfb     = -1.0434      u0      = 0.039        ua      = 0.6e-09      ub      = 1.3e-018   
+uc      = -0e-011      vsat    = 250000       a0      = 0            ags     = 0e-020     
+a1      = 0            a2      = 0.999999999  b0      = 0e-020       b1      = 0          
+keta    = 0.00         dwg     = 0            dwb     = 0            pclm    = 0.001
+pdiblc1 = 0            pdiblc2 = 0.000000001  pdiblcb = 0.000        drout   = 0.45       
+pvag    = 0e-020       delta   = 0.0189       pscbe1  = 0.00e+000    pscbe2  = 1e-10     
+fprout  = 0.0          pdits   = 0.12         pditsd  = 0.00         pditsl  = 0   
+rsh     = 0            rdsw    = 200          rsw     = 100          rdw     = 100        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 0          
+prwb    = 0e-011       wr      = 1            alpha0  = 0.074        alpha1  = 0.005      
+beta0   = 30           agidl   = 0.0002       bgidl   = 2.1e+009     cgidl   = 0.0002     
+egidl   = 0.8          

+aigbacc = 0.012        bigbacc = 0.0028       cigbacc = 0.002
+nigbacc = 1e-8         aigbinv = 0.014        bigbinv = 0.004        cigbinv = 0.004
+eigbinv = 1.1          nigbinv = 1e-8         aigc    = 0.012        bigc    = 0.0028
+cigc    = 0.002        aigsd   = 0.012        bigsd   = 0.0028       cigsd   = 0.002
+nigc    = 1e-8         poxedge = 1            pigcd   = 1            ntox    = 1

+xrcrg1  = 12           xrcrg2  = 5          
+cgso    = 2.1e-010     cgdo    = 2.1e-010     cgbo    = 2.56e-011    cgdl    = 2.495e-10     
+cgsl    = 2.495e-10    ckappas = 0.01         ckappad = 0.01         acde    = 1          
+moin    = 15           noff    = 0.9          voffcv  = 0.02       

+kt1     = -0.37        kt1l    = 0.0           kt2     = -0.042        ute     = -1.5
+ua1     = 1e-009    ub1     = -3.5e-019    uc1     = 0    prt     = 0
+at      = 53000

+fnoimod = 1            tnoimod = 0          

+jss     = 0.0001       jsws    = 1e-011       jswgs   = 1e-010       njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 1            cjs     = 0.0005       mjs     = 0.5          pbsws   = 1          
+cjsws   = 5e-010       mjsws   = 0.33         pbswgs  = 1            cjswgs  = 3e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.005        tcj     = 0.001      
+tpbsw   = 0.005        tcjsw   = 0.001        tpbswg  = 0.005        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          

+dmcg    = 0e-006       dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0.0e-008     xgw     = 0e-007       xgl     = 0e-008     

+rshg    = 0.4          gbmin   = 1e-010       rbpb    = 5            rbpd    = 15         
+rbps    = 15           rbdb    = 15           rbsb    = 15           ngcon   = 1 


* PTM 32nm PMOS
 
.model  pmos  pmos  level = 54

+version = 4.0          binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 1          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0          

+tnom    = 27           toxe    = 1.5e-009     toxp    = 8e-010       toxm    = 1.5e-009   
+dtox    = 7e-010       epsrox  = 3.9          wint    = 0e-009       lint    = 8.5e-009   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 1.5e-009   

+vth0    = -0.41174     k1      = 0.5          k2      = 0.0          k3      = 0          
+k3b     = 0            w0      = 2.5e-006     dvt0    = 1            dvt1    = 0.95        
+dvt2    = 0            dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 0.36         minv    = 0.0          voffl   = 0            dvtp0   = 0e-008     
+dvtp1   = 0.0          lpe0    = 0e-008       lpeb    = 0e-010       xj      = 1.5e-008     
+ngate   = 5e+020       ndep    = 3.5e+018     nsd     = 2e+020       phin    = 0          
+cdsc    = 0.05         cdscb   = 0            cdscd   = 0.02         cit     = 0          
+voff    = -0.155       nfactor = 1.6          eta0    = 0.035         etab    = 0          
+vfb     = 1.0642       u0      = 0.011337     ua      = 8e-010       ub      = 2.5e-018     
+uc      = 0            vsat    = 76130        a0      = 0            ags     = 0e-020     
+a1      = 0            a2      = 0.999        b0      = -1e-020      b1      = 0          
+keta    = 0.0          dwg     = 0            dwb     = 0            pclm    = 0.001       
+pdiblc1 = 0.0          pdiblc2 = 0.0000001    pdiblcb = 0            drout   = 0.45       
+pvag    = 0e-020       delta   = 0.04         pscbe1  = 0e+00        pscbe2  = 1e-010  
+fprout  = 0.0          pdits   = 0.15         pditsd  = 0.0          pditsl  = 0   
+rsh     = 0            rdsw    = 300          rsw     = 150          rdw     = 150        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 0
+prwb    = 0            wr      = 1            alpha0  = 0.074        alpha1  = 0.005      
+beta0   = 30           agidl   = 0.0002       bgidl   = 2.1e+009     cgidl   = 0.0002     
+egidl   = 0.8          

+aigbacc = 0.012        bigbacc = 0.0028       cigbacc = 0.002
+nigbacc = 1            aigbinv = 0.014        bigbinv = 0.004        cigbinv = 0.004
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.69         bigc    = 0.0012
+cigc    = 0.0008       aigsd   = 0.0087       bigsd   = 0.0012       cigsd   = 0.0008
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1

+xrcrg1  = 12           xrcrg2  = 5          
+cgso    = 2.1e-010     cgdo    = 2.1e-010     cgbo    = 2.56e-011    cgdl    = 1e-014     
+cgsl    = 1e-014       ckappas = 0.5          ckappad = 0.5          acde    = 1          
+moin    = 15           noff    = 0.9          voffcv  = 0.02       

+kt1     = -0.34        kt1l    = 0            kt2     = -0.052        ute     = -1.5
+ua1     = -1e-009    ub1     = 2e-018    uc1     = 0    prt     = 0
+at      = 33000

+fnoimod = 1            tnoimod = 0          

+jss     = 0.0001       jsws    = 1e-011       jswgs   = 1e-010       njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 1            cjs     = 0.0005       mjs     = 0.5          pbsws   = 1          
+cjsws   = 5e-010       mjsws   = 0.33         pbswgs  = 1            cjswgs  = 3e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.005        tcj     = 0.001      
+tpbsw   = 0.005        tcjsw   = 0.001        tpbswg  = 0.005        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          

+dmcg    = 0e-006       dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0e-008     xgw     = 0e-007       xgl     = 0e-008     

+rshg    = 0.4          gbmin   = 1e-010       rbpb    = 5            rbpd    = 15         
+rbps    = 15           rbdb    = 15           rbsb    = 15           ngcon   = 1 

.end